library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.ALL;

entity mux is 
port(
    RegDst_in   : in STD_LOGIC;
    Branch_in   : in STD_LOGIC;
    MemRead_in  : in STD_LOGIC;
    MemtoReg_in : in STD_LOGIC;
    MemWrite_in : in STD_LOGIC;
    ALUSrc_in   : in STD_LOGIC;
    RegWrite_in : in STD_LOGIC;
    Jump_in     : in STD_LOGIC;
    ALUOp_in    : in STD_LOGIC_VECTOR(1 downto 0);
    sel         : in std_logic;

    RegDst_out  : out STD_LOGIC;
    Branch_out  : out STD_LOGIC;
    MemRead_out : out STD_LOGIC;
    MemtoReg_out    : out STD_LOGIC;
    MemWrite_out    : out STD_LOGIC;
    ALUSrc_out  : out STD_LOGIC;
    RegWrite_out    : out STD_LOGIC;
    Jump_out    : out STD_LOGIC;
    ALUOp_out   : out STD_LOGIC_VECTOR(1 downto 0)
);
end mux;

architecture arch of mux is
begin
	process(RegDst_in,Branch_in,MemRead_in,MemtoReg_in,MemWrite_in,ALUSrc_in,RegWrite_in,Jump_in,ALUOp_in,sel)
	begin
		if(sel = '0') then
			RegDst_out <= RegDst_in;
			Branch_out <= Branch_in;
			MemRead_out <= MemRead_in;
			MemtoReg_out <= MemtoReg_in;
			MemWrite_out <= MemWrite_in;
			ALUSrc_out <= ALUSrc_in;
			RegWrite_out <= RegWrite_in;
			Jump_out <= Jump_in;
			ALUOp_out <= ALUOp_in;
		else
			RegDst_out <= '0';
			Branch_out <= '0';
			MemRead_out <= '0';
			MemtoReg_out <= '0';
			MemWrite_out <= '0';
			ALUSrc_out <= '0';
			RegWrite_out <= '0';
			Jump_out <= '0';
			ALUOp_out <= "00";
		end if;
	end process;
end arch;

--worked with Ruoxi



			
